<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-11.8559,-19.2127,129.627,-89.145</PageViewport>
<gate>
<ID>28</ID>
<type>AE_SMALL_INVERTER</type>
<position>58,-27</position>
<input>
<ID>IN_0</ID>5 </input>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_TOGGLE</type>
<position>52,-27</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>32</ID>
<type>GA_LED</type>
<position>62.5,-27</position>
<input>
<ID>N_in0</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>57,-24.5</position>
<gparam>LABEL_TEXT NOT Gate</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>52,-33</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_TOGGLE</type>
<position>52,-37</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_AND2</type>
<position>58,-35</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>GA_LED</type>
<position>62.5,-35</position>
<input>
<ID>N_in0</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>AA_LABEL</type>
<position>57,-30</position>
<gparam>LABEL_TEXT AND Gate</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>57,-39</position>
<gparam>LABEL_TEXT OR Gate</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>AE_OR2</type>
<position>58,-44</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_TOGGLE</type>
<position>52,-42</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_TOGGLE</type>
<position>52,-46</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>52</ID>
<type>GA_LED</type>
<position>62.5,-44</position>
<input>
<ID>N_in0</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>AA_LABEL</type>
<position>57,-48.5</position>
<gparam>LABEL_TEXT NAND Gate</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>AA_TOGGLE</type>
<position>52,-52</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_TOGGLE</type>
<position>52,-56</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>59</ID>
<type>BA_NAND2</type>
<position>58,-54</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>61</ID>
<type>GA_LED</type>
<position>62.5,-54</position>
<input>
<ID>N_in0</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>AA_LABEL</type>
<position>57,-58.5</position>
<gparam>LABEL_TEXT NOR Gate</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>AA_TOGGLE</type>
<position>52,-62</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>66</ID>
<type>AA_TOGGLE</type>
<position>52,-66</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>68</ID>
<type>BE_NOR2</type>
<position>58,-64</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>18 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>70</ID>
<type>GA_LED</type>
<position>62.5,-64</position>
<input>
<ID>N_in0</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>71</ID>
<type>AA_LABEL</type>
<position>57,-68.5</position>
<gparam>LABEL_TEXT XOR Gate</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>73</ID>
<type>AA_TOGGLE</type>
<position>52,-72</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>75</ID>
<type>AA_TOGGLE</type>
<position>52,-76</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>77</ID>
<type>AI_XOR2</type>
<position>58,-74</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>79</ID>
<type>GA_LED</type>
<position>62.5,-74</position>
<input>
<ID>N_in0</ID>21 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>80</ID>
<type>AA_LABEL</type>
<position>57,-78.5</position>
<gparam>LABEL_TEXT XNOR Gate</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>AA_TOGGLE</type>
<position>52,-82</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_TOGGLE</type>
<position>52,-86</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>86</ID>
<type>GA_LED</type>
<position>62.5,-84</position>
<input>
<ID>N_in0</ID>24 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>AO_XNOR2</type>
<position>58,-84</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>89</ID>
<type>AA_LABEL</type>
<position>67,-27</position>
<gparam>LABEL_TEXT Y = A'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>AA_LABEL</type>
<position>67.5,-34.5</position>
<gparam>LABEL_TEXT Y = A.B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>AA_LABEL</type>
<position>68,-43.5</position>
<gparam>LABEL_TEXT Y = A+B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>AA_LABEL</type>
<position>68.5,-53.5</position>
<gparam>LABEL_TEXT Y = (A.B)'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>93</ID>
<type>AA_LABEL</type>
<position>68.5,-63.5</position>
<gparam>LABEL_TEXT Y = (A+B)'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>94</ID>
<type>AA_LABEL</type>
<position>72,-73.5</position>
<gparam>LABEL_TEXT Y = ((A.B')+(A'.B))</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>95</ID>
<type>AA_LABEL</type>
<position>72,-83.5</position>
<gparam>LABEL_TEXT Y = ((A.B)+(A'.B'))</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,-27,56,-27</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<intersection>56 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>56,-27,56,-27</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>-27 1</intersection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-27,61.5,-27</points>
<connection>
<GID>32</GID>
<name>N_in0</name></connection>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-34,54.5,-33</points>
<intersection>-34 1</intersection>
<intersection>-33 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-34,55,-34</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54,-33,54.5,-33</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-37,54.5,-36</points>
<intersection>-37 2</intersection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-36,55,-36</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54,-37,54.5,-37</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61,-35,61.5,-35</points>
<connection>
<GID>40</GID>
<name>OUT</name></connection>
<connection>
<GID>42</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-43,54.5,-42</points>
<intersection>-43 1</intersection>
<intersection>-42 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-43,55,-43</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54,-42,54.5,-42</points>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-46,54.5,-45</points>
<intersection>-46 2</intersection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-45,55,-45</points>
<connection>
<GID>46</GID>
<name>IN_1</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54,-46,54.5,-46</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61,-44,61.5,-44</points>
<connection>
<GID>46</GID>
<name>OUT</name></connection>
<connection>
<GID>52</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-53,54.5,-52</points>
<intersection>-53 1</intersection>
<intersection>-52 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-53,55,-53</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54,-52,54.5,-52</points>
<connection>
<GID>55</GID>
<name>OUT_0</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-56,54.5,-55</points>
<intersection>-56 2</intersection>
<intersection>-55 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-55,55,-55</points>
<connection>
<GID>59</GID>
<name>IN_1</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54,-56,54.5,-56</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61,-54,61.5,-54</points>
<connection>
<GID>59</GID>
<name>OUT</name></connection>
<connection>
<GID>61</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61,-64,61.5,-64</points>
<connection>
<GID>68</GID>
<name>OUT</name></connection>
<connection>
<GID>70</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-63,54.5,-62</points>
<intersection>-63 1</intersection>
<intersection>-62 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-63,55,-63</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54,-62,54.5,-62</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-66,54.5,-65</points>
<intersection>-66 2</intersection>
<intersection>-65 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-65,55,-65</points>
<connection>
<GID>68</GID>
<name>IN_1</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54,-66,54.5,-66</points>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-73,54.5,-72</points>
<intersection>-73 1</intersection>
<intersection>-72 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-73,55,-73</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54,-72,54.5,-72</points>
<connection>
<GID>73</GID>
<name>OUT_0</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-76,54.5,-75</points>
<intersection>-76 2</intersection>
<intersection>-75 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-75,55,-75</points>
<connection>
<GID>77</GID>
<name>IN_1</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54,-76,54.5,-76</points>
<connection>
<GID>75</GID>
<name>OUT_0</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61,-74,61.5,-74</points>
<connection>
<GID>77</GID>
<name>OUT</name></connection>
<connection>
<GID>79</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-83,54.5,-82</points>
<intersection>-83 1</intersection>
<intersection>-82 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-83,55,-83</points>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54,-82,54.5,-82</points>
<connection>
<GID>82</GID>
<name>OUT_0</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-86,54.5,-85</points>
<intersection>-86 2</intersection>
<intersection>-85 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-85,55,-85</points>
<connection>
<GID>88</GID>
<name>IN_1</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54,-86,54.5,-86</points>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61,-84,61.5,-84</points>
<connection>
<GID>88</GID>
<name>OUT</name></connection>
<connection>
<GID>86</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-831.914,20.2652,-545.686,-121.212</PageViewport>
<gate>
<ID>103</ID>
<type>AA_LABEL</type>
<position>-691.5,-10.5</position>
<gparam>LABEL_TEXT NOT Gate (Y=A')</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>105</ID>
<type>AA_TOGGLE</type>
<position>-699,-14</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>107</ID>
<type>BA_NAND2</type>
<position>-691.5,-14</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>27 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>111</ID>
<type>GA_LED</type>
<position>-686,-14</position>
<input>
<ID>N_in0</ID>28 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>113</ID>
<type>AA_TOGGLE</type>
<position>-699,-19</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>115</ID>
<type>BE_NOR2</type>
<position>-691.5,-19</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>117</ID>
<type>GA_LED</type>
<position>-686,-19</position>
<input>
<ID>N_in0</ID>30 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>AA_LABEL</type>
<position>-693,-24</position>
<gparam>LABEL_TEXT AND Gate (Y=(A.B))</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>120</ID>
<type>AA_TOGGLE</type>
<position>-703,-27</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>122</ID>
<type>AA_TOGGLE</type>
<position>-703,-31</position>
<output>
<ID>OUT_0</ID>33 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>124</ID>
<type>BA_NAND2</type>
<position>-696,-29</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>126</ID>
<type>BA_NAND2</type>
<position>-689,-29</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>128</ID>
<type>GA_LED</type>
<position>-684,-29</position>
<input>
<ID>N_in0</ID>35 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>130</ID>
<type>AA_TOGGLE</type>
<position>-703,-36</position>
<output>
<ID>OUT_0</ID>38 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>132</ID>
<type>AA_TOGGLE</type>
<position>-703,-41</position>
<output>
<ID>OUT_0</ID>39 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>136</ID>
<type>BE_NOR2</type>
<position>-696,-36</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>138</ID>
<type>BE_NOR2</type>
<position>-696,-41</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>39 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>140</ID>
<type>BE_NOR2</type>
<position>-689,-38.5</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>41 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>142</ID>
<type>GA_LED</type>
<position>-684,-38.5</position>
<input>
<ID>N_in0</ID>42 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>143</ID>
<type>AA_LABEL</type>
<position>-693,-45</position>
<gparam>LABEL_TEXT OR Gate (Y=(A+B))</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>145</ID>
<type>AA_TOGGLE</type>
<position>-703,-50</position>
<output>
<ID>OUT_0</ID>43 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>147</ID>
<type>AA_TOGGLE</type>
<position>-703,-56</position>
<output>
<ID>OUT_0</ID>45 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>149</ID>
<type>BA_NAND2</type>
<position>-696,-50</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>43 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>151</ID>
<type>BA_NAND2</type>
<position>-696,-56</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>45 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>153</ID>
<type>BA_NAND2</type>
<position>-688,-53</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>48 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>155</ID>
<type>GA_LED</type>
<position>-683,-53</position>
<input>
<ID>N_in0</ID>49 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>157</ID>
<type>AA_TOGGLE</type>
<position>-703,-61</position>
<output>
<ID>OUT_0</ID>50 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>159</ID>
<type>BE_NOR2</type>
<position>-696,-63</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>51 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>161</ID>
<type>AA_TOGGLE</type>
<position>-703,-65</position>
<output>
<ID>OUT_0</ID>51 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>163</ID>
<type>BE_NOR2</type>
<position>-689,-63</position>
<input>
<ID>IN_0</ID>52 </input>
<input>
<ID>IN_1</ID>52 </input>
<output>
<ID>OUT</ID>53 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>165</ID>
<type>GA_LED</type>
<position>-683,-63</position>
<input>
<ID>N_in0</ID>53 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>166</ID>
<type>AA_LABEL</type>
<position>-692.5,-68.5</position>
<gparam>LABEL_TEXT NAND Gate (Y = (A.B)')</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>169</ID>
<type>AA_TOGGLE</type>
<position>-705,-74</position>
<output>
<ID>OUT_0</ID>54 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>170</ID>
<type>AA_TOGGLE</type>
<position>-705,-79</position>
<output>
<ID>OUT_0</ID>55 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>171</ID>
<type>BE_NOR2</type>
<position>-698,-74</position>
<input>
<ID>IN_0</ID>54 </input>
<input>
<ID>IN_1</ID>54 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>172</ID>
<type>BE_NOR2</type>
<position>-698,-79</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>55 </input>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>173</ID>
<type>BE_NOR2</type>
<position>-691,-76.5</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>57 </input>
<output>
<ID>OUT</ID>59 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>176</ID>
<type>BE_NOR2</type>
<position>-684,-76.5</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>59 </input>
<output>
<ID>OUT</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>178</ID>
<type>GA_LED</type>
<position>-680,-76.5</position>
<input>
<ID>N_in0</ID>60 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>179</ID>
<type>AA_LABEL</type>
<position>-691.5,-83</position>
<gparam>LABEL_TEXT NOR Gate (Y = (A+B)')</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>180</ID>
<type>AA_TOGGLE</type>
<position>-705,-88</position>
<output>
<ID>OUT_0</ID>61 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>181</ID>
<type>AA_TOGGLE</type>
<position>-705,-94</position>
<output>
<ID>OUT_0</ID>62 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>182</ID>
<type>BA_NAND2</type>
<position>-698,-88</position>
<input>
<ID>IN_0</ID>61 </input>
<input>
<ID>IN_1</ID>61 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>183</ID>
<type>BA_NAND2</type>
<position>-698,-94</position>
<input>
<ID>IN_0</ID>62 </input>
<input>
<ID>IN_1</ID>62 </input>
<output>
<ID>OUT</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>184</ID>
<type>BA_NAND2</type>
<position>-690,-91</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>64 </input>
<output>
<ID>OUT</ID>66 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>187</ID>
<type>BA_NAND2</type>
<position>-683,-91</position>
<input>
<ID>IN_0</ID>66 </input>
<input>
<ID>IN_1</ID>66 </input>
<output>
<ID>OUT</ID>67 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>189</ID>
<type>GA_LED</type>
<position>-679,-91</position>
<input>
<ID>N_in0</ID>67 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>190</ID>
<type>AA_LABEL</type>
<position>-690.5,-98.5</position>
<gparam>LABEL_TEXT XOR Gate (Y = ((A.B')+(A'.B)))</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-694.5,-15,-694.5,-13</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<connection>
<GID>107</GID>
<name>IN_1</name></connection>
<intersection>-14 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-697,-14,-694.5,-14</points>
<connection>
<GID>105</GID>
<name>OUT_0</name></connection>
<intersection>-694.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-688.5,-14,-687,-14</points>
<connection>
<GID>111</GID>
<name>N_in0</name></connection>
<connection>
<GID>107</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-694.5,-20,-694.5,-18</points>
<connection>
<GID>115</GID>
<name>IN_1</name></connection>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-697,-19,-694.5,-19</points>
<connection>
<GID>113</GID>
<name>OUT_0</name></connection>
<intersection>-694.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-688.5,-19,-687,-19</points>
<connection>
<GID>117</GID>
<name>N_in0</name></connection>
<connection>
<GID>115</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-700,-28,-700,-27</points>
<intersection>-28 3</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-701,-27,-700,-27</points>
<connection>
<GID>120</GID>
<name>OUT_0</name></connection>
<intersection>-700 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-700,-28,-699,-28</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>-700 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-700,-31,-700,-30</points>
<intersection>-31 2</intersection>
<intersection>-30 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-701,-31,-700,-31</points>
<connection>
<GID>122</GID>
<name>OUT_0</name></connection>
<intersection>-700 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-700,-30,-699,-30</points>
<connection>
<GID>124</GID>
<name>IN_1</name></connection>
<intersection>-700 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-692,-30,-692,-28</points>
<connection>
<GID>126</GID>
<name>IN_1</name></connection>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-693,-29,-692,-29</points>
<connection>
<GID>124</GID>
<name>OUT</name></connection>
<intersection>-692 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-686,-29,-685,-29</points>
<connection>
<GID>126</GID>
<name>OUT</name></connection>
<connection>
<GID>128</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-699,-37,-699,-35</points>
<connection>
<GID>136</GID>
<name>IN_1</name></connection>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-701,-36,-699,-36</points>
<connection>
<GID>130</GID>
<name>OUT_0</name></connection>
<intersection>-699 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-699,-42,-699,-40</points>
<connection>
<GID>138</GID>
<name>IN_1</name></connection>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>-41 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-701,-41,-699,-41</points>
<connection>
<GID>132</GID>
<name>OUT_0</name></connection>
<intersection>-699 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-692.5,-37.5,-692.5,-36</points>
<intersection>-37.5 1</intersection>
<intersection>-36 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-692.5,-37.5,-692,-37.5</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>-692.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-693,-36,-692.5,-36</points>
<connection>
<GID>136</GID>
<name>OUT</name></connection>
<intersection>-692.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-692.5,-41,-692.5,-39.5</points>
<intersection>-41 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-692.5,-39.5,-692,-39.5</points>
<connection>
<GID>140</GID>
<name>IN_1</name></connection>
<intersection>-692.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-693,-41,-692.5,-41</points>
<connection>
<GID>138</GID>
<name>OUT</name></connection>
<intersection>-692.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-686,-38.5,-685,-38.5</points>
<connection>
<GID>142</GID>
<name>N_in0</name></connection>
<connection>
<GID>140</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-699,-51,-699,-49</points>
<connection>
<GID>149</GID>
<name>IN_1</name></connection>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<intersection>-50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-701,-50,-699,-50</points>
<connection>
<GID>145</GID>
<name>OUT_0</name></connection>
<intersection>-699 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-699,-57,-699,-55</points>
<connection>
<GID>151</GID>
<name>IN_1</name></connection>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-701,-56,-699,-56</points>
<connection>
<GID>147</GID>
<name>OUT_0</name></connection>
<intersection>-699 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-692,-52,-692,-50</points>
<intersection>-52 1</intersection>
<intersection>-50 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-692,-52,-691,-52</points>
<connection>
<GID>153</GID>
<name>IN_0</name></connection>
<intersection>-692 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-693,-50,-692,-50</points>
<connection>
<GID>149</GID>
<name>OUT</name></connection>
<intersection>-692 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-692,-56,-692,-54</points>
<intersection>-56 2</intersection>
<intersection>-54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-692,-54,-691,-54</points>
<connection>
<GID>153</GID>
<name>IN_1</name></connection>
<intersection>-692 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-693,-56,-692,-56</points>
<connection>
<GID>151</GID>
<name>OUT</name></connection>
<intersection>-692 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-685,-53,-684,-53</points>
<connection>
<GID>155</GID>
<name>N_in0</name></connection>
<connection>
<GID>153</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-701,-61,-699,-61</points>
<connection>
<GID>157</GID>
<name>OUT_0</name></connection>
<intersection>-699 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-699,-62,-699,-61</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>-61 1</intersection></vsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-699,-65,-699,-64</points>
<connection>
<GID>159</GID>
<name>IN_1</name></connection>
<intersection>-65 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-701,-65,-699,-65</points>
<connection>
<GID>161</GID>
<name>OUT_0</name></connection>
<intersection>-699 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-692,-64,-692,-62</points>
<connection>
<GID>163</GID>
<name>IN_1</name></connection>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-693,-63,-692,-63</points>
<connection>
<GID>159</GID>
<name>OUT</name></connection>
<intersection>-692 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-686,-63,-684,-63</points>
<connection>
<GID>163</GID>
<name>OUT</name></connection>
<connection>
<GID>165</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-701,-75,-701,-73</points>
<connection>
<GID>171</GID>
<name>IN_1</name></connection>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>-74 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-703,-74,-701,-74</points>
<connection>
<GID>169</GID>
<name>OUT_0</name></connection>
<intersection>-701 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-701,-80,-701,-78</points>
<connection>
<GID>172</GID>
<name>IN_1</name></connection>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-703,-79,-701,-79</points>
<connection>
<GID>170</GID>
<name>OUT_0</name></connection>
<intersection>-701 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-694.5,-75.5,-694.5,-74</points>
<intersection>-75.5 1</intersection>
<intersection>-74 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-694.5,-75.5,-694,-75.5</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<intersection>-694.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-695,-74,-694.5,-74</points>
<connection>
<GID>171</GID>
<name>OUT</name></connection>
<intersection>-694.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-694.5,-79,-694.5,-77.5</points>
<intersection>-79 2</intersection>
<intersection>-77.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-694.5,-77.5,-694,-77.5</points>
<connection>
<GID>173</GID>
<name>IN_1</name></connection>
<intersection>-694.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-695,-79,-694.5,-79</points>
<connection>
<GID>172</GID>
<name>OUT</name></connection>
<intersection>-694.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-687,-77.5,-687,-75.5</points>
<connection>
<GID>176</GID>
<name>IN_1</name></connection>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>-76.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-688,-76.5,-687,-76.5</points>
<connection>
<GID>173</GID>
<name>OUT</name></connection>
<intersection>-687 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-681,-76.5,-681,-76.5</points>
<connection>
<GID>176</GID>
<name>OUT</name></connection>
<connection>
<GID>178</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-701,-89,-701,-87</points>
<connection>
<GID>182</GID>
<name>IN_1</name></connection>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>-88 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-703,-88,-701,-88</points>
<connection>
<GID>180</GID>
<name>OUT_0</name></connection>
<intersection>-701 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-701,-95,-701,-93</points>
<connection>
<GID>183</GID>
<name>IN_1</name></connection>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>-94 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-703,-94,-701,-94</points>
<connection>
<GID>181</GID>
<name>OUT_0</name></connection>
<intersection>-701 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-694,-90,-694,-88</points>
<intersection>-90 1</intersection>
<intersection>-88 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-694,-90,-693,-90</points>
<connection>
<GID>184</GID>
<name>IN_0</name></connection>
<intersection>-694 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-695,-88,-694,-88</points>
<connection>
<GID>182</GID>
<name>OUT</name></connection>
<intersection>-694 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-694,-94,-694,-92</points>
<intersection>-94 2</intersection>
<intersection>-92 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-694,-92,-693,-92</points>
<connection>
<GID>184</GID>
<name>IN_1</name></connection>
<intersection>-694 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-695,-94,-694,-94</points>
<connection>
<GID>183</GID>
<name>OUT</name></connection>
<intersection>-694 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-686,-92,-686,-90</points>
<connection>
<GID>187</GID>
<name>IN_1</name></connection>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<intersection>-91 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-687,-91,-686,-91</points>
<connection>
<GID>184</GID>
<name>OUT</name></connection>
<intersection>-686 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-680,-91,-680,-91</points>
<connection>
<GID>187</GID>
<name>OUT</name></connection>
<connection>
<GID>189</GID>
<name>N_in0</name></connection></vsegment></shape></wire></page 1>
<page 2>
<PageViewport>34,-19.7622,88.4,-46.651</PageViewport>
<gate>
<ID>194</ID>
<type>AA_TOGGLE</type>
<position>53,-29</position>
<output>
<ID>OUT_0</ID>68 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>196</ID>
<type>AA_TOGGLE</type>
<position>53,-33</position>
<output>
<ID>OUT_0</ID>69 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>198</ID>
<type>AI_XOR2</type>
<position>60,-31</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>69 </input>
<output>
<ID>OUT</ID>70 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>200</ID>
<type>AA_AND2</type>
<position>60,-36</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>69 </input>
<output>
<ID>OUT</ID>71 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>202</ID>
<type>GA_LED</type>
<position>64,-31</position>
<input>
<ID>N_in0</ID>70 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>204</ID>
<type>GA_LED</type>
<position>64,-36</position>
<input>
<ID>N_in0</ID>71 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>192</ID>
<type>AA_LABEL</type>
<position>58,-25.5</position>
<gparam>LABEL_TEXT Half Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>68</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-29,57,-29</points>
<connection>
<GID>194</GID>
<name>OUT_0</name></connection>
<intersection>56.5 3</intersection>
<intersection>57 6</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>56.5,-35,56.5,-29</points>
<intersection>-35 5</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>56.5,-35,57,-35</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<intersection>56.5 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>57,-30,57,-29</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<intersection>-29 1</intersection></vsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-37,56,-32</points>
<intersection>-37 3</intersection>
<intersection>-33 2</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-32,57,-32</points>
<connection>
<GID>198</GID>
<name>IN_1</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55,-33,56,-33</points>
<connection>
<GID>196</GID>
<name>OUT_0</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>56,-37,57,-37</points>
<connection>
<GID>200</GID>
<name>IN_1</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-31,63,-31</points>
<connection>
<GID>198</GID>
<name>OUT</name></connection>
<connection>
<GID>202</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-36,63,-36</points>
<connection>
<GID>200</GID>
<name>OUT</name></connection>
<connection>
<GID>204</GID>
<name>N_in0</name></connection></vsegment></shape></wire></page 2>
<page 3>
<PageViewport>26.775,-18.275,95.625,-52.3063</PageViewport>
<gate>
<ID>206</ID>
<type>AA_TOGGLE</type>
<position>50,-26</position>
<output>
<ID>OUT_0</ID>73 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>208</ID>
<type>AA_LABEL</type>
<position>56.5,-21.5</position>
<gparam>LABEL_TEXT Full Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>210</ID>
<type>AA_TOGGLE</type>
<position>50,-29</position>
<output>
<ID>OUT_0</ID>74 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>212</ID>
<type>AA_TOGGLE</type>
<position>50,-32</position>
<output>
<ID>OUT_0</ID>75 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>216</ID>
<type>AI_XOR3</type>
<position>60,-29</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>74 </input>
<input>
<ID>IN_2</ID>75 </input>
<output>
<ID>OUT</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>218</ID>
<type>GA_LED</type>
<position>64,-29</position>
<input>
<ID>N_in0</ID>76 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>220</ID>
<type>AA_AND2</type>
<position>60,-36</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>222</ID>
<type>AA_AND2</type>
<position>60,-41</position>
<input>
<ID>IN_0</ID>74 </input>
<input>
<ID>IN_1</ID>75 </input>
<output>
<ID>OUT</ID>82 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>224</ID>
<type>AA_AND2</type>
<position>60,-46</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>73 </input>
<output>
<ID>OUT</ID>83 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>230</ID>
<type>AE_OR3</type>
<position>67.5,-41</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>82 </input>
<input>
<ID>IN_2</ID>83 </input>
<output>
<ID>OUT</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>232</ID>
<type>GA_LED</type>
<position>71.5,-41</position>
<input>
<ID>N_in0</ID>84 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-27,55,-26</points>
<intersection>-27 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-27,57,-27</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<intersection>54 3</intersection>
<intersection>55 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52,-26,55,-26</points>
<connection>
<GID>206</GID>
<name>OUT_0</name></connection>
<intersection>55 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>54,-47,54,-27</points>
<intersection>-47 4</intersection>
<intersection>-45 6</intersection>
<intersection>-35 7</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>54,-47,57,-47</points>
<connection>
<GID>224</GID>
<name>IN_1</name></connection>
<intersection>54 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>54,-45,57,-45</points>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<intersection>54 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>54,-35,57,-35</points>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<intersection>54 3</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52,-29,57,-29</points>
<connection>
<GID>216</GID>
<name>IN_1</name></connection>
<connection>
<GID>210</GID>
<name>OUT_0</name></connection>
<intersection>55 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>55,-40,55,-29</points>
<intersection>-40 4</intersection>
<intersection>-37 5</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>55,-40,57,-40</points>
<connection>
<GID>222</GID>
<name>IN_0</name></connection>
<intersection>55 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>55,-37,57,-37</points>
<connection>
<GID>220</GID>
<name>IN_1</name></connection>
<intersection>55 3</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-42,56,-31</points>
<intersection>-42 3</intersection>
<intersection>-32 2</intersection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-31,57,-31</points>
<connection>
<GID>216</GID>
<name>IN_2</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52,-32,56,-32</points>
<connection>
<GID>212</GID>
<name>OUT_0</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>56,-42,57,-42</points>
<connection>
<GID>222</GID>
<name>IN_1</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-29,63,-29</points>
<connection>
<GID>216</GID>
<name>OUT</name></connection>
<connection>
<GID>218</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-39,63.5,-36</points>
<intersection>-39 1</intersection>
<intersection>-36 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-39,64.5,-39</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63,-36,63.5,-36</points>
<connection>
<GID>220</GID>
<name>OUT</name></connection>
<intersection>63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>63,-41,64.5,-41</points>
<connection>
<GID>230</GID>
<name>IN_1</name></connection>
<connection>
<GID>222</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-46,63.5,-43</points>
<intersection>-46 2</intersection>
<intersection>-43 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-43,64.5,-43</points>
<connection>
<GID>230</GID>
<name>IN_2</name></connection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63,-46,63.5,-46</points>
<connection>
<GID>224</GID>
<name>OUT</name></connection>
<intersection>63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-41,70.5,-41</points>
<connection>
<GID>230</GID>
<name>OUT</name></connection>
<connection>
<GID>232</GID>
<name>N_in0</name></connection></vsegment></shape></wire></page 3>
<page 4>
<PageViewport>24.4385,-8.45547,97.9615,-44.7965</PageViewport>
<gate>
<ID>234</ID>
<type>AA_FULLADDER_1BIT</type>
<position>47,-27</position>
<input>
<ID>IN_0</ID>92 </input>
<input>
<ID>IN_B_0</ID>93 </input>
<output>
<ID>OUT_0</ID>94 </output>
<input>
<ID>carry_in</ID>103 </input>
<output>
<ID>carry_out</ID>106 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>236</ID>
<type>AA_FULLADDER_1BIT</type>
<position>57,-27</position>
<input>
<ID>IN_0</ID>90 </input>
<input>
<ID>IN_B_0</ID>91 </input>
<output>
<ID>OUT_0</ID>95 </output>
<input>
<ID>carry_in</ID>104 </input>
<output>
<ID>carry_out</ID>103 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>238</ID>
<type>AA_FULLADDER_1BIT</type>
<position>67,-27</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_B_0</ID>89 </input>
<output>
<ID>OUT_0</ID>96 </output>
<input>
<ID>carry_in</ID>98 </input>
<output>
<ID>carry_out</ID>104 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>240</ID>
<type>AA_FULLADDER_1BIT</type>
<position>77,-27</position>
<input>
<ID>IN_0</ID>108 </input>
<input>
<ID>IN_B_0</ID>87 </input>
<output>
<ID>OUT_0</ID>97 </output>
<input>
<ID>carry_in</ID>107 </input>
<output>
<ID>carry_out</ID>98 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>242</ID>
<type>AA_LABEL</type>
<position>61,-16.5</position>
<gparam>LABEL_TEXT An Adder which can Add 2 singal digits</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>244</ID>
<type>FF_GND</type>
<position>82,-27</position>
<output>
<ID>OUT_0</ID>107 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>246</ID>
<type>AA_TOGGLE</type>
<position>79,-20</position>
<output>
<ID>OUT_0</ID>108 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>247</ID>
<type>AA_TOGGLE</type>
<position>75,-20</position>
<output>
<ID>OUT_0</ID>87 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>248</ID>
<type>AA_TOGGLE</type>
<position>69,-20</position>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>249</ID>
<type>AA_TOGGLE</type>
<position>65,-20</position>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>250</ID>
<type>AA_TOGGLE</type>
<position>59,-20</position>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>251</ID>
<type>AA_TOGGLE</type>
<position>55,-20</position>
<output>
<ID>OUT_0</ID>91 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>252</ID>
<type>AA_TOGGLE</type>
<position>49,-20</position>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>253</ID>
<type>AA_TOGGLE</type>
<position>45,-20</position>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>255</ID>
<type>GA_LED</type>
<position>47,-31</position>
<input>
<ID>N_in3</ID>94 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>257</ID>
<type>GA_LED</type>
<position>57,-31</position>
<input>
<ID>N_in3</ID>95 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>259</ID>
<type>GA_LED</type>
<position>67,-31</position>
<input>
<ID>N_in3</ID>96 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>261</ID>
<type>GA_LED</type>
<position>77,-31</position>
<input>
<ID>N_in3</ID>97 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>267</ID>
<type>GA_LED</type>
<position>42,-27</position>
<input>
<ID>N_in1</ID>106 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>269</ID>
<type>AA_LABEL</type>
<position>60.5,-33.5</position>
<gparam>LABEL_TEXT 4-bit Parallel Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-23,75,-22</points>
<connection>
<GID>247</GID>
<name>OUT_0</name></connection>
<intersection>-23 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>76,-24,76,-23</points>
<connection>
<GID>240</GID>
<name>IN_B_0</name></connection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>75,-23,76,-23</points>
<intersection>75 0</intersection>
<intersection>76 1</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-23,69,-22</points>
<connection>
<GID>248</GID>
<name>OUT_0</name></connection>
<intersection>-23 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>68,-24,68,-23</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>68,-23,69,-23</points>
<intersection>68 1</intersection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-23,65,-22</points>
<connection>
<GID>249</GID>
<name>OUT_0</name></connection>
<intersection>-23 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>66,-24,66,-23</points>
<connection>
<GID>238</GID>
<name>IN_B_0</name></connection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>65,-23,66,-23</points>
<intersection>65 0</intersection>
<intersection>66 1</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59,-23,59,-22</points>
<connection>
<GID>250</GID>
<name>OUT_0</name></connection>
<intersection>-23 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>58,-24,58,-23</points>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>58,-23,59,-23</points>
<intersection>58 1</intersection>
<intersection>59 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-23,55,-22</points>
<connection>
<GID>251</GID>
<name>OUT_0</name></connection>
<intersection>-23 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>56,-24,56,-23</points>
<connection>
<GID>236</GID>
<name>IN_B_0</name></connection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>55,-23,56,-23</points>
<intersection>55 0</intersection>
<intersection>56 1</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-23,49,-22</points>
<connection>
<GID>252</GID>
<name>OUT_0</name></connection>
<intersection>-23 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>48,-24,48,-23</points>
<connection>
<GID>234</GID>
<name>IN_0</name></connection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>48,-23,49,-23</points>
<intersection>48 1</intersection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-23,45,-22</points>
<connection>
<GID>253</GID>
<name>OUT_0</name></connection>
<intersection>-23 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>46,-24,46,-23</points>
<connection>
<GID>234</GID>
<name>IN_B_0</name></connection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>45,-23,46,-23</points>
<intersection>45 0</intersection>
<intersection>46 1</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-30,47,-30</points>
<connection>
<GID>234</GID>
<name>OUT_0</name></connection>
<connection>
<GID>255</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-30,57,-30</points>
<connection>
<GID>236</GID>
<name>OUT_0</name></connection>
<connection>
<GID>257</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-30,67,-30</points>
<connection>
<GID>238</GID>
<name>OUT_0</name></connection>
<connection>
<GID>259</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,-30,77,-30</points>
<connection>
<GID>240</GID>
<name>OUT_0</name></connection>
<connection>
<GID>261</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-27,73,-27</points>
<connection>
<GID>240</GID>
<name>carry_out</name></connection>
<connection>
<GID>238</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51,-27,53,-27</points>
<connection>
<GID>236</GID>
<name>carry_out</name></connection>
<connection>
<GID>234</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61,-27,63,-27</points>
<connection>
<GID>238</GID>
<name>carry_out</name></connection>
<connection>
<GID>236</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-27,43,-27</points>
<connection>
<GID>234</GID>
<name>carry_out</name></connection>
<connection>
<GID>267</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-27,81,-27</points>
<connection>
<GID>240</GID>
<name>carry_in</name></connection>
<connection>
<GID>244</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-24,78,-23</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<intersection>-23 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>79,-23,79,-22</points>
<connection>
<GID>246</GID>
<name>OUT_0</name></connection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>78,-23,79,-23</points>
<intersection>78 0</intersection>
<intersection>79 1</intersection></hsegment></shape></wire></page 4>
<page 5>
<PageViewport>10.2375,7.6375,102.037,-37.7375</PageViewport>
<gate>
<ID>271</ID>
<type>AE_FULLADDER_4BIT</type>
<position>53,-22.5</position>
<input>
<ID>IN_0</ID>134 </input>
<input>
<ID>IN_1</ID>135 </input>
<input>
<ID>IN_2</ID>136 </input>
<input>
<ID>IN_3</ID>137 </input>
<input>
<ID>IN_B_0</ID>133 </input>
<input>
<ID>IN_B_1</ID>132 </input>
<input>
<ID>IN_B_2</ID>131 </input>
<input>
<ID>IN_B_3</ID>130 </input>
<output>
<ID>OUT_0</ID>138 </output>
<output>
<ID>OUT_1</ID>139 </output>
<output>
<ID>OUT_2</ID>140 </output>
<output>
<ID>OUT_3</ID>141 </output>
<input>
<ID>carry_in</ID>113 </input>
<output>
<ID>carry_out</ID>143 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>275</ID>
<type>FF_GND</type>
<position>62.5,-21.5</position>
<output>
<ID>OUT_0</ID>113 </output>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>277</ID>
<type>DD_KEYPAD_HEX</type>
<position>41,-12.5</position>
<output>
<ID>OUT_0</ID>134 </output>
<output>
<ID>OUT_1</ID>135 </output>
<output>
<ID>OUT_2</ID>136 </output>
<output>
<ID>OUT_3</ID>137 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 8</lparam></gate>
<gate>
<ID>279</ID>
<type>DD_KEYPAD_HEX</type>
<position>41,0.5</position>
<output>
<ID>OUT_0</ID>133 </output>
<output>
<ID>OUT_1</ID>132 </output>
<output>
<ID>OUT_2</ID>131 </output>
<output>
<ID>OUT_3</ID>130 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 8</lparam></gate>
<gate>
<ID>283</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>65,-30.5</position>
<input>
<ID>IN_0</ID>138 </input>
<input>
<ID>IN_1</ID>139 </input>
<input>
<ID>IN_2</ID>140 </input>
<input>
<ID>IN_3</ID>141 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>287</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>41.5,-30.5</position>
<input>
<ID>IN_0</ID>143 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>289</ID>
<type>AA_LABEL</type>
<position>77.5,-5.5</position>
<gparam>LABEL_TEXT An Adder which can Add 2 singal digits</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>291</ID>
<type>AA_LABEL</type>
<position>77,-9</position>
<gparam>LABEL_TEXT 4-Bit Full Adder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>113</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61,-21.5,61.5,-21.5</points>
<connection>
<GID>275</GID>
<name>OUT_0</name></connection>
<connection>
<GID>271</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-18.5,55,3.5</points>
<connection>
<GID>271</GID>
<name>IN_B_3</name></connection>
<intersection>3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,3.5,55,3.5</points>
<connection>
<GID>279</GID>
<name>OUT_3</name></connection>
<intersection>55 0</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-18.5,56,1.5</points>
<connection>
<GID>271</GID>
<name>IN_B_2</name></connection>
<intersection>1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,1.5,56,1.5</points>
<connection>
<GID>279</GID>
<name>OUT_2</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-18.5,57,-0.5</points>
<connection>
<GID>271</GID>
<name>IN_B_1</name></connection>
<intersection>-0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-0.5,57,-0.5</points>
<connection>
<GID>279</GID>
<name>OUT_1</name></connection>
<intersection>57 0</intersection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,-18.5,58,-2.5</points>
<connection>
<GID>271</GID>
<name>IN_B_0</name></connection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-2.5,58,-2.5</points>
<connection>
<GID>279</GID>
<name>OUT_0</name></connection>
<intersection>58 0</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-18.5,51,-15.5</points>
<connection>
<GID>271</GID>
<name>IN_0</name></connection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-15.5,51,-15.5</points>
<connection>
<GID>277</GID>
<name>OUT_0</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-18.5,50,-13.5</points>
<connection>
<GID>271</GID>
<name>IN_1</name></connection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-13.5,50,-13.5</points>
<connection>
<GID>277</GID>
<name>OUT_1</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-18.5,49,-11.5</points>
<connection>
<GID>271</GID>
<name>IN_2</name></connection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-11.5,49,-11.5</points>
<connection>
<GID>277</GID>
<name>OUT_2</name></connection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-18.5,48,-9.5</points>
<connection>
<GID>271</GID>
<name>IN_3</name></connection>
<intersection>-9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-9.5,48,-9.5</points>
<connection>
<GID>277</GID>
<name>OUT_3</name></connection>
<intersection>48 0</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-31.5,54.5,-26.5</points>
<connection>
<GID>271</GID>
<name>OUT_0</name></connection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-31.5,62,-31.5</points>
<connection>
<GID>283</GID>
<name>IN_0</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-30.5,53.5,-26.5</points>
<connection>
<GID>271</GID>
<name>OUT_1</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53.5,-30.5,62,-30.5</points>
<connection>
<GID>283</GID>
<name>IN_1</name></connection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-29.5,52.5,-26.5</points>
<connection>
<GID>271</GID>
<name>OUT_2</name></connection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52.5,-29.5,62,-29.5</points>
<connection>
<GID>283</GID>
<name>IN_2</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-28.5,51.5,-26.5</points>
<connection>
<GID>271</GID>
<name>OUT_3</name></connection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51.5,-28.5,62,-28.5</points>
<connection>
<GID>283</GID>
<name>IN_3</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-31.5,35,-21.5</points>
<intersection>-31.5 1</intersection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-31.5,38.5,-31.5</points>
<connection>
<GID>287</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,-21.5,45,-21.5</points>
<connection>
<GID>271</GID>
<name>carry_out</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire></page 5>
<page 6>
<PageViewport>20.025,-9.8375,88.875,-43.8688</PageViewport>
<gate>
<ID>293</ID>
<type>AI_XOR2</type>
<position>52,-21</position>
<input>
<ID>IN_0</ID>144 </input>
<input>
<ID>IN_1</ID>145 </input>
<output>
<ID>OUT</ID>147 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>295</ID>
<type>AA_TOGGLE</type>
<position>39.5,-20</position>
<output>
<ID>OUT_0</ID>144 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>297</ID>
<type>AA_TOGGLE</type>
<position>39.5,-25</position>
<output>
<ID>OUT_0</ID>145 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>299</ID>
<type>AA_AND2</type>
<position>52,-32.5</position>
<input>
<ID>IN_0</ID>149 </input>
<input>
<ID>IN_1</ID>145 </input>
<output>
<ID>OUT</ID>148 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>303</ID>
<type>GA_LED</type>
<position>56,-21</position>
<input>
<ID>N_in0</ID>147 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>305</ID>
<type>GA_LED</type>
<position>56,-32.5</position>
<input>
<ID>N_in0</ID>148 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>307</ID>
<type>AE_SMALL_INVERTER</type>
<position>45.5,-28.5</position>
<input>
<ID>IN_0</ID>144 </input>
<output>
<ID>OUT_0</ID>149 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>309</ID>
<type>AA_LABEL</type>
<position>62,-20.5</position>
<gparam>LABEL_TEXT Difference</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>310</ID>
<type>AA_LABEL</type>
<position>60.5,-32</position>
<gparam>LABEL_TEXT Borrow</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>311</ID>
<type>AA_LABEL</type>
<position>53.5,-15.5</position>
<gparam>LABEL_TEXT Half Subtractor</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>144</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41.5,-20,49,-20</points>
<connection>
<GID>293</GID>
<name>IN_0</name></connection>
<connection>
<GID>295</GID>
<name>OUT_0</name></connection>
<intersection>45.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>45.5,-26.5,45.5,-20</points>
<connection>
<GID>307</GID>
<name>IN_0</name></connection>
<intersection>-20 1</intersection></vsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-33.5,48,-22</points>
<intersection>-33.5 3</intersection>
<intersection>-25 2</intersection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,-22,49,-22</points>
<connection>
<GID>293</GID>
<name>IN_1</name></connection>
<intersection>48 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41.5,-25,48,-25</points>
<connection>
<GID>297</GID>
<name>OUT_0</name></connection>
<intersection>48 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>48,-33.5,49,-33.5</points>
<connection>
<GID>299</GID>
<name>IN_1</name></connection>
<intersection>48 0</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-21,55,-21</points>
<connection>
<GID>293</GID>
<name>OUT</name></connection>
<connection>
<GID>303</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-32.5,55,-32.5</points>
<connection>
<GID>305</GID>
<name>N_in0</name></connection>
<connection>
<GID>299</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-31.5,45.5,-30.5</points>
<connection>
<GID>307</GID>
<name>OUT_0</name></connection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45.5,-31.5,49,-31.5</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<intersection>45.5 0</intersection></hsegment></shape></wire></page 6>
<page 7>
<PageViewport>20.025,-16.5875,88.875,-50.6188</PageViewport>
<gate>
<ID>313</ID>
<type>AA_LABEL</type>
<position>52,-18</position>
<gparam>LABEL_TEXT Full Subtractor</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>315</ID>
<type>AI_XOR3</type>
<position>53,-25</position>
<input>
<ID>IN_0</ID>150 </input>
<input>
<ID>IN_1</ID>151 </input>
<input>
<ID>IN_2</ID>152 </input>
<output>
<ID>OUT</ID>157 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>317</ID>
<type>AA_TOGGLE</type>
<position>40,-22</position>
<output>
<ID>OUT_0</ID>150 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>319</ID>
<type>AA_TOGGLE</type>
<position>40,-25</position>
<output>
<ID>OUT_0</ID>151 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>321</ID>
<type>AA_TOGGLE</type>
<position>40,-28</position>
<output>
<ID>OUT_0</ID>152 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>323</ID>
<type>AE_SMALL_INVERTER</type>
<position>44.5,-31.5</position>
<input>
<ID>IN_0</ID>150 </input>
<output>
<ID>OUT_0</ID>153 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>325</ID>
<type>AA_AND2</type>
<position>53,-35</position>
<input>
<ID>IN_0</ID>153 </input>
<input>
<ID>IN_1</ID>152 </input>
<output>
<ID>OUT</ID>154 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>327</ID>
<type>AA_AND2</type>
<position>53,-40</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>152 </input>
<output>
<ID>OUT</ID>155 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>329</ID>
<type>AA_AND2</type>
<position>53,-45</position>
<input>
<ID>IN_0</ID>153 </input>
<input>
<ID>IN_1</ID>151 </input>
<output>
<ID>OUT</ID>156 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>331</ID>
<type>AE_OR3</type>
<position>60,-40</position>
<input>
<ID>IN_0</ID>154 </input>
<input>
<ID>IN_1</ID>155 </input>
<input>
<ID>IN_2</ID>156 </input>
<output>
<ID>OUT</ID>158 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>333</ID>
<type>GA_LED</type>
<position>57,-25</position>
<input>
<ID>N_in0</ID>157 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>335</ID>
<type>GA_LED</type>
<position>64,-40</position>
<input>
<ID>N_in0</ID>158 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>336</ID>
<type>AA_LABEL</type>
<position>63,-25</position>
<gparam>LABEL_TEXT Difference</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>337</ID>
<type>AA_LABEL</type>
<position>68.5,-40</position>
<gparam>LABEL_TEXT Borrow</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-29.5,44.5,-22</points>
<connection>
<GID>323</GID>
<name>IN_0</name></connection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42,-22,49.5,-22</points>
<connection>
<GID>317</GID>
<name>OUT_0</name></connection>
<intersection>44.5 0</intersection>
<intersection>49.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>49.5,-23,49.5,-22</points>
<intersection>-23 4</intersection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>49.5,-23,50,-23</points>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<intersection>49.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42,-25,50,-25</points>
<connection>
<GID>319</GID>
<name>OUT_0</name></connection>
<connection>
<GID>315</GID>
<name>IN_1</name></connection>
<intersection>46 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>46,-46,46,-25</points>
<intersection>-46 12</intersection>
<intersection>-39 10</intersection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>46,-39,50,-39</points>
<connection>
<GID>327</GID>
<name>IN_0</name></connection>
<intersection>46 9</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>46,-46,50,-46</points>
<connection>
<GID>329</GID>
<name>IN_1</name></connection>
<intersection>46 9</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-41,43,-27</points>
<intersection>-41 7</intersection>
<intersection>-36 3</intersection>
<intersection>-28 2</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43,-27,50,-27</points>
<connection>
<GID>315</GID>
<name>IN_2</name></connection>
<intersection>43 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>42,-28,43,-28</points>
<connection>
<GID>321</GID>
<name>OUT_0</name></connection>
<intersection>43 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>43,-36,50,-36</points>
<connection>
<GID>325</GID>
<name>IN_1</name></connection>
<intersection>43 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>43,-41,50,-41</points>
<connection>
<GID>327</GID>
<name>IN_1</name></connection>
<intersection>43 0</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44.5,-34,50,-34</points>
<connection>
<GID>325</GID>
<name>IN_0</name></connection>
<intersection>44.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>44.5,-44,44.5,-33.5</points>
<connection>
<GID>323</GID>
<name>OUT_0</name></connection>
<intersection>-44 7</intersection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>44.5,-44,50,-44</points>
<connection>
<GID>329</GID>
<name>IN_0</name></connection>
<intersection>44.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-38,56.5,-35</points>
<intersection>-38 1</intersection>
<intersection>-35 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56.5,-38,57,-38</points>
<connection>
<GID>331</GID>
<name>IN_0</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56,-35,56.5,-35</points>
<connection>
<GID>325</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>56,-40,57,-40</points>
<connection>
<GID>331</GID>
<name>IN_1</name></connection>
<connection>
<GID>327</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-45,56.5,-42</points>
<intersection>-45 2</intersection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56.5,-42,57,-42</points>
<connection>
<GID>331</GID>
<name>IN_2</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56,-45,56.5,-45</points>
<connection>
<GID>329</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-25,56,-25</points>
<connection>
<GID>333</GID>
<name>N_in0</name></connection>
<connection>
<GID>315</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-40,63,-40</points>
<connection>
<GID>335</GID>
<name>N_in0</name></connection>
<connection>
<GID>331</GID>
<name>OUT</name></connection></vsegment></shape></wire></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>