<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-137.907,443.043,201.429,275.316</PageViewport>
<gate>
<ID>2</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>39,368.5</position>
<output>
<ID>A_equal_B</ID>2 </output>
<output>
<ID>A_greater_B</ID>1 </output>
<output>
<ID>A_less_B</ID>3 </output>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>9 </input>
<input>
<ID>IN_2</ID>10 </input>
<input>
<ID>IN_3</ID>11 </input>
<input>
<ID>IN_B_0</ID>4 </input>
<input>
<ID>IN_B_1</ID>5 </input>
<input>
<ID>IN_B_2</ID>6 </input>
<input>
<ID>IN_B_3</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>4</ID>
<type>GA_LED</type>
<position>29,372</position>
<input>
<ID>N_in1</ID>1 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>GA_LED</type>
<position>29,368.5</position>
<input>
<ID>N_in1</ID>2 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>29,365</position>
<input>
<ID>N_in1</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>DD_KEYPAD_HEX</type>
<position>27,391.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<output>
<ID>OUT_1</ID>5 </output>
<output>
<ID>OUT_2</ID>6 </output>
<output>
<ID>OUT_3</ID>7 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>12</ID>
<type>DD_KEYPAD_HEX</type>
<position>27,379.5</position>
<output>
<ID>OUT_0</ID>8 </output>
<output>
<ID>OUT_1</ID>9 </output>
<output>
<ID>OUT_2</ID>10 </output>
<output>
<ID>OUT_3</ID>11 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>35,401.5</position>
<gparam>LABEL_TEXT 4-bit comparator</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,370.5,30.5,372</points>
<intersection>370.5 1</intersection>
<intersection>372 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,370.5,31,370.5</points>
<connection>
<GID>2</GID>
<name>A_greater_B</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30,372,30.5,372</points>
<connection>
<GID>4</GID>
<name>N_in1</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30,368.5,31,368.5</points>
<connection>
<GID>6</GID>
<name>N_in1</name></connection>
<connection>
<GID>2</GID>
<name>A_equal_B</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,365,30.5,366.5</points>
<intersection>365 2</intersection>
<intersection>366.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,366.5,31,366.5</points>
<connection>
<GID>2</GID>
<name>A_less_B</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30,365,30.5,365</points>
<connection>
<GID>8</GID>
<name>N_in1</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,372.5,44,388.5</points>
<connection>
<GID>2</GID>
<name>IN_B_0</name></connection>
<intersection>388.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,388.5,44,388.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>44 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,372.5,43,390.5</points>
<connection>
<GID>2</GID>
<name>IN_B_1</name></connection>
<intersection>390.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,390.5,43,390.5</points>
<connection>
<GID>10</GID>
<name>OUT_1</name></connection>
<intersection>43 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,372.5,42,392.5</points>
<connection>
<GID>2</GID>
<name>IN_B_2</name></connection>
<intersection>392.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,392.5,42,392.5</points>
<connection>
<GID>10</GID>
<name>OUT_2</name></connection>
<intersection>42 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,372.5,41,394.5</points>
<connection>
<GID>2</GID>
<name>IN_B_3</name></connection>
<intersection>394.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,394.5,41,394.5</points>
<connection>
<GID>10</GID>
<name>OUT_3</name></connection>
<intersection>41 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,372.5,37,376.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>376.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,376.5,37,376.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,372.5,36,378.5</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>378.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,378.5,36,378.5</points>
<connection>
<GID>12</GID>
<name>OUT_1</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,372.5,35,380.5</points>
<connection>
<GID>2</GID>
<name>IN_2</name></connection>
<intersection>380.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,380.5,35,380.5</points>
<connection>
<GID>12</GID>
<name>OUT_2</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,372.5,34,382.5</points>
<connection>
<GID>2</GID>
<name>IN_3</name></connection>
<intersection>382.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,382.5,34,382.5</points>
<connection>
<GID>12</GID>
<name>OUT_3</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-0.704223,50.7685,296.289,-96.0294</PageViewport>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>139,2</position>
<gparam>LABEL_TEXT Draw waveform for various flipflop</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AE_DFF_LOW</type>
<position>147,-8</position>
<input>
<ID>IN_0</ID>16 </input>
<output>
<ID>OUTINV_0</ID>13 </output>
<output>
<ID>OUT_0</ID>12 </output>
<input>
<ID>clock</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>20</ID>
<type>BE_JKFF_LOW</type>
<position>147,-18.5</position>
<input>
<ID>J</ID>17 </input>
<input>
<ID>K</ID>18 </input>
<output>
<ID>Q</ID>14 </output>
<input>
<ID>clock</ID>21 </input>
<output>
<ID>nQ</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>22</ID>
<type>GA_LED</type>
<position>151,-6</position>
<input>
<ID>N_in0</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>GA_LED</type>
<position>151,-9</position>
<input>
<ID>N_in0</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>GA_LED</type>
<position>151,-16.5</position>
<input>
<ID>N_in0</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>GA_LED</type>
<position>151,-20.5</position>
<input>
<ID>N_in0</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>121,-7.5</position>
<gparam>LABEL_TEXT D-FF</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>121,-17.5</position>
<gparam>LABEL_TEXT JK-FF</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_TOGGLE</type>
<position>139,-6</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>139,-15</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_TOGGLE</type>
<position>139,-22</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>40</ID>
<type>BB_CLOCK</type>
<position>133,-10.5</position>
<output>
<ID>CLK</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>42</ID>
<type>BB_CLOCK</type>
<position>133,-18.5</position>
<output>
<ID>CLK</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>44</ID>
<type>BE_JKFF_LOW</type>
<position>147,-33</position>
<input>
<ID>J</ID>23 </input>
<input>
<ID>K</ID>23 </input>
<output>
<ID>Q</ID>25 </output>
<input>
<ID>clock</ID>24 </input>
<output>
<ID>nQ</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_TOGGLE</type>
<position>139,-31</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>50</ID>
<type>BB_CLOCK</type>
<position>133,-33</position>
<output>
<ID>CLK</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>52</ID>
<type>GA_LED</type>
<position>151,-31</position>
<input>
<ID>N_in0</ID>25 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>GA_LED</type>
<position>151,-35</position>
<input>
<ID>N_in0</ID>26 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>AA_LABEL</type>
<position>121,-32</position>
<gparam>LABEL_TEXT T-FF</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,-6,150,-6</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<connection>
<GID>22</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,-9,150,-9</points>
<connection>
<GID>18</GID>
<name>OUTINV_0</name></connection>
<connection>
<GID>24</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,-16.5,150,-16.5</points>
<connection>
<GID>20</GID>
<name>Q</name></connection>
<connection>
<GID>26</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,-20.5,150,-20.5</points>
<connection>
<GID>20</GID>
<name>nQ</name></connection>
<connection>
<GID>28</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>141,-6,144,-6</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144,-16.5,144,-15</points>
<connection>
<GID>20</GID>
<name>J</name></connection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141,-15,144,-15</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>144 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144,-22,144,-20.5</points>
<connection>
<GID>20</GID>
<name>K</name></connection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141,-22,144,-22</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<intersection>144 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140.5,-10.5,140.5,-9</points>
<intersection>-10.5 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>140.5,-9,144,-9</points>
<connection>
<GID>18</GID>
<name>clock</name></connection>
<intersection>140.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>137,-10.5,140.5,-10.5</points>
<connection>
<GID>40</GID>
<name>CLK</name></connection>
<intersection>140.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>137,-18.5,144,-18.5</points>
<connection>
<GID>20</GID>
<name>clock</name></connection>
<connection>
<GID>42</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>141,-31,144,-31</points>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<connection>
<GID>44</GID>
<name>J</name></connection>
<intersection>142.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>142.5,-35,142.5,-31</points>
<intersection>-35 3</intersection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>142.5,-35,144,-35</points>
<connection>
<GID>44</GID>
<name>K</name></connection>
<intersection>142.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>137,-33,144,-33</points>
<connection>
<GID>44</GID>
<name>clock</name></connection>
<connection>
<GID>50</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,-31,150,-31</points>
<connection>
<GID>44</GID>
<name>Q</name></connection>
<connection>
<GID>52</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,-35,150,-35</points>
<connection>
<GID>44</GID>
<name>nQ</name></connection>
<connection>
<GID>54</GID>
<name>N_in0</name></connection></vsegment></shape></wire></page 1>
<page 2>
<PageViewport>73.0937,12.8776,240.15,-69.6954</PageViewport>
<gate>
<ID>57</ID>
<type>BE_JKFF_LOW</type>
<position>159.5,-29.5</position>
<input>
<ID>J</ID>31 </input>
<input>
<ID>K</ID>33 </input>
<output>
<ID>Q</ID>34 </output>
<input>
<ID>clock</ID>32 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>59</ID>
<type>AA_TOGGLE</type>
<position>146,-24</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>61</ID>
<type>DE_TO</type>
<position>150,-24</position>
<input>
<ID>IN_0</ID>27 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID J</lparam></gate>
<gate>
<ID>67</ID>
<type>BB_CLOCK</type>
<position>139.5,-29.5</position>
<output>
<ID>CLK</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>69</ID>
<type>DE_TO</type>
<position>145.5,-29.5</position>
<input>
<ID>IN_0</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>71</ID>
<type>AA_TOGGLE</type>
<position>146,-34.5</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>73</ID>
<type>DE_TO</type>
<position>150,-34.5</position>
<input>
<ID>IN_0</ID>30 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID K</lparam></gate>
<gate>
<ID>75</ID>
<type>DA_FROM</type>
<position>154.5,-27.5</position>
<input>
<ID>IN_0</ID>31 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID J</lparam></gate>
<gate>
<ID>77</ID>
<type>DA_FROM</type>
<position>154.5,-29.5</position>
<input>
<ID>IN_0</ID>32 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>79</ID>
<type>DA_FROM</type>
<position>154.5,-31.5</position>
<input>
<ID>IN_0</ID>33 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID K</lparam></gate>
<gate>
<ID>81</ID>
<type>DE_TO</type>
<position>164.5,-27.5</position>
<input>
<ID>IN_0</ID>34 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q</lparam></gate>
<gate>
<ID>83</ID>
<type>DA_FROM</type>
<position>170,-27.5</position>
<input>
<ID>IN_0</ID>35 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q</lparam></gate>
<gate>
<ID>85</ID>
<type>GA_LED</type>
<position>173,-27.5</position>
<input>
<ID>N_in0</ID>35 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>144</ID>
<type>AA_LABEL</type>
<position>154,-15</position>
<gparam>LABEL_TEXT JK-FF Waveform</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148,-24,148,-24</points>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection>
<connection>
<GID>61</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143.5,-29.5,143.5,-29.5</points>
<connection>
<GID>67</GID>
<name>CLK</name></connection>
<connection>
<GID>69</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>148,-34.5,148,-34.5</points>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection>
<connection>
<GID>73</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-27.5,156.5,-27.5</points>
<connection>
<GID>57</GID>
<name>J</name></connection>
<connection>
<GID>75</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-29.5,156.5,-29.5</points>
<connection>
<GID>57</GID>
<name>clock</name></connection>
<connection>
<GID>77</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-31.5,156.5,-31.5</points>
<connection>
<GID>57</GID>
<name>K</name></connection>
<connection>
<GID>79</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162.5,-27.5,162.5,-27.5</points>
<connection>
<GID>57</GID>
<name>Q</name></connection>
<connection>
<GID>81</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>172,-27.5,172,-27.5</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<connection>
<GID>85</GID>
<name>N_in0</name></connection></vsegment></shape></wire></page 2>
<page 3>
<PageViewport>-17.6795,15.5943,321.657,-152.133</PageViewport>
<gate>
<ID>1</ID>
<type>BB_CLOCK</type>
<position>128.5,-47</position>
<output>
<ID>CLK</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>5</ID>
<type>GA_LED</type>
<position>182.5,-37</position>
<input>
<ID>N_in0</ID>44 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>GA_LED</type>
<position>172.5,-33</position>
<input>
<ID>N_in2</ID>28 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>GA_LED</type>
<position>158.5,-33</position>
<input>
<ID>N_in2</ID>22 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>GA_LED</type>
<position>144.5,-33</position>
<input>
<ID>N_in2</ID>19 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>BB_CLOCK</type>
<position>128.5,-68</position>
<output>
<ID>CLK</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>21</ID>
<type>GA_LED</type>
<position>182.5,-58</position>
<input>
<ID>N_in0</ID>50 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AE_DFF_LOW</type>
<position>136,-60</position>
<input>
<ID>IN_0</ID>48 </input>
<output>
<ID>OUT_0</ID>54 </output>
<input>
<ID>clock</ID>49 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>31</ID>
<type>AE_DFF_LOW</type>
<position>150,-60</position>
<input>
<ID>IN_0</ID>51 </input>
<output>
<ID>OUT_0</ID>55 </output>
<input>
<ID>clock</ID>49 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>33</ID>
<type>AE_DFF_LOW</type>
<position>163.5,-60</position>
<input>
<ID>IN_0</ID>52 </input>
<output>
<ID>OUT_0</ID>56 </output>
<input>
<ID>clock</ID>49 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>35</ID>
<type>AE_DFF_LOW</type>
<position>178.5,-60</position>
<input>
<ID>IN_0</ID>53 </input>
<output>
<ID>OUT_0</ID>50 </output>
<input>
<ID>clock</ID>49 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_TOGGLE</type>
<position>127.5,-56.5</position>
<output>
<ID>OUT_0</ID>48 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>117,-59</position>
<gparam>LABEL_TEXT PIPO</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>AA_TOGGLE</type>
<position>142.5,-52</position>
<output>
<ID>OUT_0</ID>51 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_TOGGLE</type>
<position>155.5,-52</position>
<output>
<ID>OUT_0</ID>52 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_TOGGLE</type>
<position>170,-52</position>
<output>
<ID>OUT_0</ID>53 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>53</ID>
<type>GA_LED</type>
<position>140,-58</position>
<input>
<ID>N_in0</ID>54 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>GA_LED</type>
<position>154,-58</position>
<input>
<ID>N_in0</ID>55 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>GA_LED</type>
<position>167.5,-58</position>
<input>
<ID>N_in0</ID>56 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>BB_CLOCK</type>
<position>128.5,-96.5</position>
<output>
<ID>CLK</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>64</ID>
<type>GA_LED</type>
<position>182.5,-86.5</position>
<input>
<ID>N_in0</ID>59 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>65</ID>
<type>AE_DFF_LOW</type>
<position>136,-88.5</position>
<input>
<ID>IN_0</ID>57 </input>
<output>
<ID>OUT_0</ID>67 </output>
<input>
<ID>clock</ID>58 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>66</ID>
<type>AE_DFF_LOW</type>
<position>150,-88.5</position>
<input>
<ID>IN_0</ID>69 </input>
<output>
<ID>OUT_0</ID>68 </output>
<input>
<ID>clock</ID>58 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>68</ID>
<type>AE_DFF_LOW</type>
<position>163.5,-88.5</position>
<input>
<ID>IN_0</ID>70 </input>
<output>
<ID>OUT_0</ID>71 </output>
<input>
<ID>clock</ID>58 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>70</ID>
<type>AE_DFF_LOW</type>
<position>178.5,-88.5</position>
<input>
<ID>IN_0</ID>72 </input>
<output>
<ID>OUT_0</ID>59 </output>
<input>
<ID>clock</ID>58 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>72</ID>
<type>AA_TOGGLE</type>
<position>127.5,-85</position>
<output>
<ID>OUT_0</ID>57 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_LABEL</type>
<position>117,-87.5</position>
<gparam>LABEL_TEXT PISO</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>AA_LABEL</type>
<position>153.5,-3</position>
<gparam>LABEL_TEXT Design Shift Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>AE_DFF_LOW</type>
<position>136,-15.5</position>
<input>
<ID>IN_0</ID>36 </input>
<output>
<ID>OUT_0</ID>37 </output>
<input>
<ID>clock</ID>41 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>90</ID>
<type>AA_TOGGLE</type>
<position>127.5,-77</position>
<output>
<ID>OUT_0</ID>66 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>91</ID>
<type>AE_DFF_LOW</type>
<position>148.5,-15.5</position>
<input>
<ID>IN_0</ID>37 </input>
<output>
<ID>OUT_0</ID>38 </output>
<input>
<ID>clock</ID>41 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>93</ID>
<type>AE_DFF_LOW</type>
<position>163,-15.5</position>
<input>
<ID>IN_0</ID>38 </input>
<output>
<ID>OUT_0</ID>39 </output>
<input>
<ID>clock</ID>41 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>94</ID>
<type>AA_MUX_2x1</type>
<position>142.5,-81.5</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>67 </input>
<output>
<ID>OUT</ID>69 </output>
<input>
<ID>SEL_0</ID>66 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>95</ID>
<type>AE_DFF_LOW</type>
<position>176.5,-15.5</position>
<input>
<ID>IN_0</ID>39 </input>
<output>
<ID>OUT_0</ID>40 </output>
<input>
<ID>clock</ID>41 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>97</ID>
<type>AA_TOGGLE</type>
<position>127.5,-12</position>
<output>
<ID>OUT_0</ID>36 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>98</ID>
<type>AA_MUX_2x1</type>
<position>156.5,-81.5</position>
<input>
<ID>IN_0</ID>74 </input>
<input>
<ID>IN_1</ID>68 </input>
<output>
<ID>OUT</ID>70 </output>
<input>
<ID>SEL_0</ID>66 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>99</ID>
<type>GA_LED</type>
<position>182,-12</position>
<input>
<ID>N_in0</ID>40 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>101</ID>
<type>BB_CLOCK</type>
<position>128,-25.5</position>
<output>
<ID>CLK</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>102</ID>
<type>AA_MUX_2x1</type>
<position>171,-81.5</position>
<input>
<ID>IN_0</ID>75 </input>
<input>
<ID>IN_1</ID>71 </input>
<output>
<ID>OUT</ID>72 </output>
<input>
<ID>SEL_0</ID>66 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>103</ID>
<type>AA_LABEL</type>
<position>117,-17.5</position>
<gparam>LABEL_TEXT SISO</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>105</ID>
<type>AE_DFF_LOW</type>
<position>136,-39</position>
<input>
<ID>IN_0</ID>42 </input>
<output>
<ID>OUT_0</ID>19 </output>
<input>
<ID>clock</ID>43 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>106</ID>
<type>AA_TOGGLE</type>
<position>140.5,-88</position>
<output>
<ID>OUT_0</ID>73 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>107</ID>
<type>AE_DFF_LOW</type>
<position>150,-39</position>
<input>
<ID>IN_0</ID>19 </input>
<output>
<ID>OUT_0</ID>22 </output>
<input>
<ID>clock</ID>43 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>109</ID>
<type>AE_DFF_LOW</type>
<position>163.5,-39</position>
<input>
<ID>IN_0</ID>22 </input>
<output>
<ID>OUT_0</ID>28 </output>
<input>
<ID>clock</ID>43 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>110</ID>
<type>AA_TOGGLE</type>
<position>154.5,-88</position>
<output>
<ID>OUT_0</ID>74 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>111</ID>
<type>AE_DFF_LOW</type>
<position>178.5,-39</position>
<input>
<ID>IN_0</ID>28 </input>
<output>
<ID>OUT_0</ID>44 </output>
<input>
<ID>clock</ID>43 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>113</ID>
<type>AA_TOGGLE</type>
<position>127.5,-35.5</position>
<output>
<ID>OUT_0</ID>42 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>114</ID>
<type>AA_LABEL</type>
<position>117,-38</position>
<gparam>LABEL_TEXT SIPO</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>115</ID>
<type>AA_TOGGLE</type>
<position>169,-88</position>
<output>
<ID>OUT_0</ID>75 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>116</ID>
<type>BB_CLOCK</type>
<position>129.5,-125.5</position>
<output>
<ID>CLK</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>118</ID>
<type>AE_DFF_LOW</type>
<position>137,-117.5</position>
<input>
<ID>IN_0</ID>89 </input>
<output>
<ID>OUT_0</ID>80 </output>
<input>
<ID>clock</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>119</ID>
<type>AE_DFF_LOW</type>
<position>151,-117.5</position>
<input>
<ID>IN_0</ID>82 </input>
<output>
<ID>OUT_0</ID>81 </output>
<input>
<ID>clock</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>120</ID>
<type>AE_DFF_LOW</type>
<position>164.5,-117.5</position>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>84 </output>
<input>
<ID>clock</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>121</ID>
<type>AE_DFF_LOW</type>
<position>179.5,-117.5</position>
<input>
<ID>IN_0</ID>85 </input>
<output>
<ID>OUT_0</ID>91 </output>
<input>
<ID>clock</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>123</ID>
<type>AA_LABEL</type>
<position>115,-118</position>
<gparam>LABEL_TEXT Bidirectional</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>124</ID>
<type>AA_TOGGLE</type>
<position>128.5,-106</position>
<output>
<ID>OUT_0</ID>79 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>125</ID>
<type>AA_MUX_2x1</type>
<position>143.5,-110.5</position>
<input>
<ID>IN_0</ID>84 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>82 </output>
<input>
<ID>SEL_0</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>126</ID>
<type>AA_MUX_2x1</type>
<position>157.5,-110.5</position>
<input>
<ID>IN_0</ID>91 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>83 </output>
<input>
<ID>SEL_0</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>127</ID>
<type>AA_MUX_2x1</type>
<position>172,-110.5</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>84 </input>
<output>
<ID>OUT</ID>85 </output>
<input>
<ID>SEL_0</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>130</ID>
<type>AA_TOGGLE</type>
<position>170.5,-115.5</position>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>132</ID>
<type>AA_MUX_2x1</type>
<position>131,-110.5</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>90 </input>
<output>
<ID>OUT</ID>89 </output>
<input>
<ID>SEL_0</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>134</ID>
<type>AA_TOGGLE</type>
<position>127,-109.5</position>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>136</ID>
<type>GA_LED</type>
<position>142,-116.5</position>
<input>
<ID>N_in0</ID>80 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>138</ID>
<type>GA_LED</type>
<position>156,-116.5</position>
<input>
<ID>N_in0</ID>81 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>140</ID>
<type>GA_LED</type>
<position>169.5,-118</position>
<input>
<ID>N_in0</ID>84 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>142</ID>
<type>GA_LED</type>
<position>185,-116</position>
<input>
<ID>N_in0</ID>91 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>139,-37,147,-37</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<connection>
<GID>105</GID>
<name>OUT_0</name></connection>
<intersection>144.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>144.5,-37,144.5,-34</points>
<connection>
<GID>17</GID>
<name>N_in2</name></connection>
<intersection>-37 1</intersection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>153,-37,160.5,-37</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<connection>
<GID>107</GID>
<name>OUT_0</name></connection>
<intersection>158.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>158.5,-37,158.5,-34</points>
<connection>
<GID>13</GID>
<name>N_in2</name></connection>
<intersection>-37 1</intersection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>166.5,-37,175.5,-37</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<connection>
<GID>109</GID>
<name>OUT_0</name></connection>
<intersection>172.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>172.5,-37,172.5,-34</points>
<connection>
<GID>9</GID>
<name>N_in2</name></connection>
<intersection>-37 1</intersection></vsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131,-13.5,131,-12</points>
<intersection>-13.5 1</intersection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131,-13.5,133,-13.5</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>131 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>129.5,-12,131,-12</points>
<connection>
<GID>97</GID>
<name>OUT_0</name></connection>
<intersection>131 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>139,-13.5,145.5,-13.5</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<connection>
<GID>89</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151.5,-13.5,160,-13.5</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<connection>
<GID>91</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>166,-13.5,173.5,-13.5</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<connection>
<GID>93</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179.5,-13.5,179.5,-12</points>
<connection>
<GID>95</GID>
<name>OUT_0</name></connection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>179.5,-12,181,-12</points>
<connection>
<GID>99</GID>
<name>N_in0</name></connection>
<intersection>179.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,-25.5,132,-21</points>
<connection>
<GID>101</GID>
<name>CLK</name></connection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132,-21,173.5,-21</points>
<intersection>132 0</intersection>
<intersection>133 10</intersection>
<intersection>145.5 9</intersection>
<intersection>160 8</intersection>
<intersection>173.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>173.5,-21,173.5,-16.5</points>
<connection>
<GID>95</GID>
<name>clock</name></connection>
<intersection>-21 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>160,-21,160,-16.5</points>
<connection>
<GID>93</GID>
<name>clock</name></connection>
<intersection>-21 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>145.5,-21,145.5,-16.5</points>
<connection>
<GID>91</GID>
<name>clock</name></connection>
<intersection>-21 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>133,-21,133,-16.5</points>
<connection>
<GID>89</GID>
<name>clock</name></connection>
<intersection>-21 1</intersection></vsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-37,133,-35.5</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129.5,-35.5,133,-35.5</points>
<connection>
<GID>113</GID>
<name>OUT_0</name></connection>
<intersection>133 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-47,133,-40</points>
<connection>
<GID>105</GID>
<name>clock</name></connection>
<intersection>-47 2</intersection>
<intersection>-44.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>132.5,-47,133,-47</points>
<connection>
<GID>1</GID>
<name>CLK</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>133,-44.5,175.5,-44.5</points>
<intersection>133 0</intersection>
<intersection>147 8</intersection>
<intersection>160.5 7</intersection>
<intersection>175.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>175.5,-44.5,175.5,-40</points>
<connection>
<GID>111</GID>
<name>clock</name></connection>
<intersection>-44.5 3</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>160.5,-44.5,160.5,-40</points>
<connection>
<GID>109</GID>
<name>clock</name></connection>
<intersection>-44.5 3</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>147,-44.5,147,-40</points>
<connection>
<GID>107</GID>
<name>clock</name></connection>
<intersection>-44.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181.5,-37,181.5,-37</points>
<connection>
<GID>111</GID>
<name>OUT_0</name></connection>
<connection>
<GID>5</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-58,133,-56.5</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>-56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129.5,-56.5,133,-56.5</points>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection>
<intersection>133 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-68,133,-61</points>
<connection>
<GID>29</GID>
<name>clock</name></connection>
<intersection>-68 2</intersection>
<intersection>-65.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>132.5,-68,133,-68</points>
<connection>
<GID>19</GID>
<name>CLK</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>133,-65.5,175.5,-65.5</points>
<intersection>133 0</intersection>
<intersection>147 8</intersection>
<intersection>160.5 7</intersection>
<intersection>175.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>175.5,-65.5,175.5,-61</points>
<connection>
<GID>35</GID>
<name>clock</name></connection>
<intersection>-65.5 3</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>160.5,-65.5,160.5,-61</points>
<connection>
<GID>33</GID>
<name>clock</name></connection>
<intersection>-65.5 3</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>147,-65.5,147,-61</points>
<connection>
<GID>31</GID>
<name>clock</name></connection>
<intersection>-65.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181.5,-58,181.5,-58</points>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection>
<connection>
<GID>21</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145.5,-58,145.5,-52</points>
<intersection>-58 1</intersection>
<intersection>-52 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145.5,-58,147,-58</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>145.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>144.5,-52,145.5,-52</points>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection>
<intersection>145.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159,-58,159,-52</points>
<intersection>-58 1</intersection>
<intersection>-52 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>159,-58,160.5,-58</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>159 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157.5,-52,159,-52</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>159 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173.5,-58,173.5,-52</points>
<intersection>-58 1</intersection>
<intersection>-52 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>173.5,-58,175.5,-58</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>173.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>172,-52,173.5,-52</points>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection>
<intersection>173.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,-58,139,-58</points>
<connection>
<GID>53</GID>
<name>N_in0</name></connection>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153,-58,153,-58</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<connection>
<GID>58</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166.5,-58,166.5,-58</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<connection>
<GID>62</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-86.5,133,-85</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>-85 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129.5,-85,133,-85</points>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<intersection>133 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-96.5,133,-89.5</points>
<connection>
<GID>65</GID>
<name>clock</name></connection>
<intersection>-96.5 2</intersection>
<intersection>-94 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>132.5,-96.5,133,-96.5</points>
<connection>
<GID>63</GID>
<name>CLK</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>133,-94,175.5,-94</points>
<intersection>133 0</intersection>
<intersection>147 8</intersection>
<intersection>160.5 7</intersection>
<intersection>175.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>175.5,-94,175.5,-89.5</points>
<connection>
<GID>70</GID>
<name>clock</name></connection>
<intersection>-94 3</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>160.5,-94,160.5,-89.5</points>
<connection>
<GID>68</GID>
<name>clock</name></connection>
<intersection>-94 3</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>147,-94,147,-89.5</points>
<connection>
<GID>66</GID>
<name>clock</name></connection>
<intersection>-94 3</intersection></vsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181.5,-86.5,181.5,-86.5</points>
<connection>
<GID>70</GID>
<name>OUT_0</name></connection>
<connection>
<GID>64</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>171,-79,171,-77</points>
<connection>
<GID>102</GID>
<name>SEL_0</name></connection>
<intersection>-77 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129.5,-77,171,-77</points>
<connection>
<GID>90</GID>
<name>OUT_0</name></connection>
<intersection>142.5 3</intersection>
<intersection>156.5 2</intersection>
<intersection>171 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>156.5,-79,156.5,-77</points>
<connection>
<GID>98</GID>
<name>SEL_0</name></connection>
<intersection>-77 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>142.5,-79,142.5,-77</points>
<connection>
<GID>94</GID>
<name>SEL_0</name></connection>
<intersection>-77 1</intersection></vsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139.5,-86.5,139.5,-80.5</points>
<intersection>-86.5 2</intersection>
<intersection>-80.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>139.5,-80.5,140.5,-80.5</points>
<connection>
<GID>94</GID>
<name>IN_1</name></connection>
<intersection>139.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>139,-86.5,139.5,-86.5</points>
<connection>
<GID>65</GID>
<name>OUT_0</name></connection>
<intersection>139.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153.5,-86.5,153.5,-80.5</points>
<intersection>-86.5 2</intersection>
<intersection>-80.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>153.5,-80.5,154.5,-80.5</points>
<connection>
<GID>98</GID>
<name>IN_1</name></connection>
<intersection>153.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>153,-86.5,153.5,-86.5</points>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection>
<intersection>153.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145.5,-86.5,145.5,-81.5</points>
<intersection>-86.5 1</intersection>
<intersection>-81.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145.5,-86.5,147,-86.5</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>145.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>144.5,-81.5,145.5,-81.5</points>
<connection>
<GID>94</GID>
<name>OUT</name></connection>
<intersection>145.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159.5,-86.5,159.5,-81.5</points>
<intersection>-86.5 1</intersection>
<intersection>-81.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>159.5,-86.5,160.5,-86.5</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>159.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>158.5,-81.5,159.5,-81.5</points>
<connection>
<GID>98</GID>
<name>OUT</name></connection>
<intersection>159.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167.5,-86.5,167.5,-80.5</points>
<intersection>-86.5 1</intersection>
<intersection>-80.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166.5,-86.5,167.5,-86.5</points>
<connection>
<GID>68</GID>
<name>OUT_0</name></connection>
<intersection>167.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>167.5,-80.5,169,-80.5</points>
<connection>
<GID>102</GID>
<name>IN_1</name></connection>
<intersection>167.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>174,-86.5,174,-81.5</points>
<intersection>-86.5 1</intersection>
<intersection>-81.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>174,-86.5,175.5,-86.5</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>174 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>173,-81.5,174,-81.5</points>
<connection>
<GID>102</GID>
<name>OUT</name></connection>
<intersection>174 0</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140.5,-86,140.5,-82.5</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<connection>
<GID>106</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>154.5,-86,154.5,-82.5</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<connection>
<GID>110</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169,-86,169,-82.5</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<connection>
<GID>115</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134,-125.5,134,-118.5</points>
<connection>
<GID>118</GID>
<name>clock</name></connection>
<intersection>-125.5 2</intersection>
<intersection>-123 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>133.5,-125.5,134,-125.5</points>
<connection>
<GID>116</GID>
<name>CLK</name></connection>
<intersection>134 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>134,-123,176.5,-123</points>
<intersection>134 0</intersection>
<intersection>148 8</intersection>
<intersection>161.5 7</intersection>
<intersection>176.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>176.5,-123,176.5,-118.5</points>
<connection>
<GID>121</GID>
<name>clock</name></connection>
<intersection>-123 3</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>161.5,-123,161.5,-118.5</points>
<connection>
<GID>120</GID>
<name>clock</name></connection>
<intersection>-123 3</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>148,-123,148,-118.5</points>
<connection>
<GID>119</GID>
<name>clock</name></connection>
<intersection>-123 3</intersection></vsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>172,-108,172,-106</points>
<connection>
<GID>127</GID>
<name>SEL_0</name></connection>
<intersection>-106 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130.5,-106,172,-106</points>
<connection>
<GID>124</GID>
<name>OUT_0</name></connection>
<intersection>131 4</intersection>
<intersection>143.5 3</intersection>
<intersection>157.5 2</intersection>
<intersection>172 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>157.5,-108,157.5,-106</points>
<connection>
<GID>126</GID>
<name>SEL_0</name></connection>
<intersection>-106 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>143.5,-108,143.5,-106</points>
<connection>
<GID>125</GID>
<name>SEL_0</name></connection>
<intersection>-106 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>131,-108,131,-106</points>
<connection>
<GID>132</GID>
<name>SEL_0</name></connection>
<intersection>-106 1</intersection></vsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140.5,-116.5,140.5,-109.5</points>
<intersection>-116.5 3</intersection>
<intersection>-115.5 2</intersection>
<intersection>-109.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>140.5,-109.5,141.5,-109.5</points>
<connection>
<GID>125</GID>
<name>IN_1</name></connection>
<intersection>140.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>140,-115.5,140.5,-115.5</points>
<connection>
<GID>118</GID>
<name>OUT_0</name></connection>
<intersection>140.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>140.5,-116.5,141,-116.5</points>
<connection>
<GID>136</GID>
<name>N_in0</name></connection>
<intersection>140.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>154.5,-110,154.5,-109.5</points>
<intersection>-110 2</intersection>
<intersection>-109.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154.5,-109.5,155.5,-109.5</points>
<connection>
<GID>126</GID>
<name>IN_1</name></connection>
<intersection>154.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>129,-110,154.5,-110</points>
<intersection>129 3</intersection>
<intersection>154 4</intersection>
<intersection>154.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>129,-111.5,129,-110</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>-110 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>154,-116.5,154,-110</points>
<connection>
<GID>119</GID>
<name>OUT_0</name></connection>
<intersection>-116.5 5</intersection>
<intersection>-110 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>154,-116.5,155,-116.5</points>
<connection>
<GID>138</GID>
<name>N_in0</name></connection>
<intersection>154 4</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146.5,-115.5,146.5,-110.5</points>
<intersection>-115.5 1</intersection>
<intersection>-110.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>146.5,-115.5,148,-115.5</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>146.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>145.5,-110.5,146.5,-110.5</points>
<connection>
<GID>125</GID>
<name>OUT</name></connection>
<intersection>146.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160.5,-115.5,160.5,-110.5</points>
<intersection>-115.5 1</intersection>
<intersection>-110.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>160.5,-115.5,161.5,-115.5</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>160.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>159.5,-110.5,160.5,-110.5</points>
<connection>
<GID>126</GID>
<name>OUT</name></connection>
<intersection>160.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168.5,-113,168.5,-109.5</points>
<intersection>-113 1</intersection>
<intersection>-109.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-113,168.5,-113</points>
<intersection>141.5 4</intersection>
<intersection>168 3</intersection>
<intersection>168.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>168.5,-109.5,170,-109.5</points>
<connection>
<GID>127</GID>
<name>IN_1</name></connection>
<intersection>168.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>168,-118,168,-113</points>
<intersection>-118 6</intersection>
<intersection>-115.5 5</intersection>
<intersection>-113 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>141.5,-113,141.5,-111.5</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>-113 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>167.5,-115.5,168,-115.5</points>
<connection>
<GID>120</GID>
<name>OUT_0</name></connection>
<intersection>168 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>168,-118,168.5,-118</points>
<connection>
<GID>140</GID>
<name>N_in0</name></connection>
<intersection>168 3</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>175,-115.5,175,-110.5</points>
<intersection>-115.5 1</intersection>
<intersection>-110.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>175,-115.5,176.5,-115.5</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>175 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>174,-110.5,175,-110.5</points>
<connection>
<GID>127</GID>
<name>OUT</name></connection>
<intersection>175 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170.5,-113.5,170.5,-111.5</points>
<connection>
<GID>130</GID>
<name>OUT_0</name></connection>
<intersection>-111.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>170,-111.5,170.5,-111.5</points>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<intersection>170.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133.5,-115.5,133.5,-110.5</points>
<intersection>-115.5 1</intersection>
<intersection>-110.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133.5,-115.5,134,-115.5</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>133.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>133,-110.5,133.5,-110.5</points>
<connection>
<GID>132</GID>
<name>OUT</name></connection>
<intersection>133.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129,-109.5,129,-109.5</points>
<connection>
<GID>132</GID>
<name>IN_1</name></connection>
<connection>
<GID>134</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169,-114,169,-113</points>
<intersection>-114 2</intersection>
<intersection>-113 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169,-113,182.5,-113</points>
<intersection>169 0</intersection>
<intersection>182.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>155.5,-114,169,-114</points>
<intersection>155.5 3</intersection>
<intersection>169 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>155.5,-114,155.5,-111.5</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<intersection>-114 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>182.5,-116,182.5,-113</points>
<connection>
<GID>121</GID>
<name>OUT_0</name></connection>
<intersection>-116 5</intersection>
<intersection>-113 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>182.5,-116,184,-116</points>
<connection>
<GID>142</GID>
<name>N_in0</name></connection>
<intersection>182.5 4</intersection></hsegment></shape></wire></page 3>
<page 4>
<PageViewport>394.381,-40.0356,496.266,-90.3954</PageViewport>
<gate>
<ID>196</ID>
<type>GA_LED</type>
<position>432.5,-24</position>
<input>
<ID>N_in2</ID>106 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>198</ID>
<type>GA_LED</type>
<position>445,-24</position>
<input>
<ID>N_in2</ID>107 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>200</ID>
<type>GA_LED</type>
<position>458.5,-24</position>
<input>
<ID>N_in2</ID>108 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>204</ID>
<type>AA_TOGGLE</type>
<position>426.5,-18</position>
<output>
<ID>OUT_0</ID>114 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>206</ID>
<type>GA_LED</type>
<position>472,-23</position>
<input>
<ID>N_in0</ID>113 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>209</ID>
<type>AA_LABEL</type>
<position>448.5,-42.5</position>
<gparam>LABEL_TEXT Johnson Counter</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>210</ID>
<type>GA_LED</type>
<position>433,-55.5</position>
<input>
<ID>N_in2</ID>116 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>211</ID>
<type>GA_LED</type>
<position>445.5,-55.5</position>
<input>
<ID>N_in2</ID>117 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>212</ID>
<type>GA_LED</type>
<position>459,-55.5</position>
<input>
<ID>N_in2</ID>118 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>214</ID>
<type>GA_LED</type>
<position>472.5,-55.5</position>
<input>
<ID>N_in2</ID>122 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>215</ID>
<type>AE_DFF_LOW</type>
<position>427,-61</position>
<input>
<ID>IN_0</ID>123 </input>
<output>
<ID>OUT_0</ID>116 </output>
<input>
<ID>clock</ID>119 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>216</ID>
<type>AE_DFF_LOW</type>
<position>439.5,-61</position>
<input>
<ID>IN_0</ID>116 </input>
<output>
<ID>OUT_0</ID>117 </output>
<input>
<ID>clock</ID>119 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>217</ID>
<type>AE_DFF_LOW</type>
<position>452,-61</position>
<input>
<ID>IN_0</ID>117 </input>
<output>
<ID>OUT_0</ID>118 </output>
<input>
<ID>clock</ID>119 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>218</ID>
<type>AE_DFF_LOW</type>
<position>466,-61</position>
<input>
<ID>IN_0</ID>118 </input>
<output>
<ID>OUTINV_0</ID>123 </output>
<output>
<ID>OUT_0</ID>122 </output>
<input>
<ID>clock</ID>119 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>219</ID>
<type>BB_CLOCK</type>
<position>420,-67.5</position>
<output>
<ID>CLK</ID>119 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>146</ID>
<type>AA_LABEL</type>
<position>446,38</position>
<gparam>LABEL_TEXT 2-Bit UP Counter</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>148</ID>
<type>BE_JKFF_LOW</type>
<position>440.5,26.5</position>
<input>
<ID>J</ID>93 </input>
<input>
<ID>K</ID>93 </input>
<output>
<ID>Q</ID>92 </output>
<input>
<ID>clock</ID>95 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>150</ID>
<type>BE_JKFF_LOW</type>
<position>458.5,26.5</position>
<input>
<ID>J</ID>92 </input>
<input>
<ID>K</ID>92 </input>
<output>
<ID>Q</ID>94 </output>
<input>
<ID>clock</ID>95 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>152</ID>
<type>AA_TOGGLE</type>
<position>430,28.5</position>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>154</ID>
<type>GA_LED</type>
<position>446,26.5</position>
<input>
<ID>N_in0</ID>92 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>156</ID>
<type>GA_LED</type>
<position>463,27</position>
<input>
<ID>N_in0</ID>94 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>158</ID>
<type>BB_CLOCK</type>
<position>430.5,20</position>
<output>
<ID>CLK</ID>95 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>159</ID>
<type>AA_LABEL</type>
<position>446.5,11.5</position>
<gparam>LABEL_TEXT 2-Bit DOWN Counter</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>160</ID>
<type>BE_JKFF_LOW</type>
<position>441.5,0.5</position>
<input>
<ID>J</ID>97 </input>
<input>
<ID>K</ID>97 </input>
<output>
<ID>Q</ID>100 </output>
<input>
<ID>clock</ID>99 </input>
<output>
<ID>nQ</ID>101 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>161</ID>
<type>BE_JKFF_LOW</type>
<position>459.5,0.5</position>
<input>
<ID>J</ID>101 </input>
<input>
<ID>K</ID>101 </input>
<output>
<ID>Q</ID>98 </output>
<input>
<ID>clock</ID>99 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>162</ID>
<type>AA_TOGGLE</type>
<position>430.5,2.5</position>
<output>
<ID>OUT_0</ID>97 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>163</ID>
<type>GA_LED</type>
<position>445.5,2.5</position>
<input>
<ID>N_in0</ID>100 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>164</ID>
<type>GA_LED</type>
<position>463.5,2.5</position>
<input>
<ID>N_in0</ID>98 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>165</ID>
<type>BB_CLOCK</type>
<position>431.5,-6</position>
<output>
<ID>CLK</ID>99 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>166</ID>
<type>AA_LABEL</type>
<position>447,-13</position>
<gparam>LABEL_TEXT RING Counter</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>174</ID>
<type>AE_DFF_LOW</type>
<position>426.5,-29.5</position>
<input>
<ID>IN_0</ID>113 </input>
<output>
<ID>OUT_0</ID>106 </output>
<input>
<ID>clock</ID>110 </input>
<input>
<ID>set</ID>114 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>176</ID>
<type>AE_DFF_LOW</type>
<position>439,-29.5</position>
<input>
<ID>IN_0</ID>106 </input>
<output>
<ID>OUT_0</ID>107 </output>
<input>
<ID>clock</ID>110 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>178</ID>
<type>AE_DFF_LOW</type>
<position>451.5,-29.5</position>
<input>
<ID>IN_0</ID>107 </input>
<output>
<ID>OUT_0</ID>108 </output>
<input>
<ID>clock</ID>110 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>180</ID>
<type>AE_DFF_LOW</type>
<position>465.5,-29.5</position>
<input>
<ID>IN_0</ID>108 </input>
<output>
<ID>OUT_0</ID>113 </output>
<input>
<ID>clock</ID>110 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>182</ID>
<type>BB_CLOCK</type>
<position>419.5,-36</position>
<output>
<ID>CLK</ID>110 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<wire>
<ID>92</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>443.5,28.5,455.5,28.5</points>
<connection>
<GID>148</GID>
<name>Q</name></connection>
<connection>
<GID>150</GID>
<name>J</name></connection>
<intersection>444.5 4</intersection>
<intersection>450 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>450,24.5,450,28.5</points>
<intersection>24.5 3</intersection>
<intersection>28.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>450,24.5,455.5,24.5</points>
<connection>
<GID>150</GID>
<name>K</name></connection>
<intersection>450 2</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>444.5,26.5,444.5,28.5</points>
<intersection>26.5 5</intersection>
<intersection>28.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>444.5,26.5,445,26.5</points>
<connection>
<GID>154</GID>
<name>N_in0</name></connection>
<intersection>444.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>432,28.5,437.5,28.5</points>
<connection>
<GID>148</GID>
<name>J</name></connection>
<connection>
<GID>152</GID>
<name>OUT_0</name></connection>
<intersection>435 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>435,24.5,435,28.5</points>
<intersection>24.5 4</intersection>
<intersection>28.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>435,24.5,437.5,24.5</points>
<connection>
<GID>148</GID>
<name>K</name></connection>
<intersection>435 3</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>461.5,27,461.5,28.5</points>
<connection>
<GID>150</GID>
<name>Q</name></connection>
<intersection>27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>461.5,27,462,27</points>
<connection>
<GID>156</GID>
<name>N_in0</name></connection>
<intersection>461.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>436,20,436,21.5</points>
<intersection>20 1</intersection>
<intersection>21.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>434.5,20,436,20</points>
<connection>
<GID>158</GID>
<name>CLK</name></connection>
<intersection>436 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>436,21.5,453.5,21.5</points>
<intersection>436 0</intersection>
<intersection>437 5</intersection>
<intersection>453.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>453.5,21.5,453.5,26.5</points>
<intersection>21.5 2</intersection>
<intersection>26.5 6</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>437,21.5,437,26.5</points>
<intersection>21.5 2</intersection>
<intersection>26.5 7</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>453.5,26.5,455.5,26.5</points>
<connection>
<GID>150</GID>
<name>clock</name></connection>
<intersection>453.5 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>437,26.5,437.5,26.5</points>
<connection>
<GID>148</GID>
<name>clock</name></connection>
<intersection>437 5</intersection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>432.5,2.5,438.5,2.5</points>
<connection>
<GID>160</GID>
<name>J</name></connection>
<connection>
<GID>162</GID>
<name>OUT_0</name></connection>
<intersection>436 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>436,-1.5,436,2.5</points>
<intersection>-1.5 4</intersection>
<intersection>2.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>436,-1.5,438.5,-1.5</points>
<connection>
<GID>160</GID>
<name>K</name></connection>
<intersection>436 3</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>462.5,2.5,462.5,2.5</points>
<connection>
<GID>161</GID>
<name>Q</name></connection>
<connection>
<GID>164</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>437,-6,437,-4.5</points>
<intersection>-6 1</intersection>
<intersection>-4.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>435.5,-6,437,-6</points>
<connection>
<GID>165</GID>
<name>CLK</name></connection>
<intersection>437 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>437,-4.5,454.5,-4.5</points>
<intersection>437 0</intersection>
<intersection>438 5</intersection>
<intersection>454.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>454.5,-4.5,454.5,0.5</points>
<intersection>-4.5 2</intersection>
<intersection>0.5 6</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>438,-4.5,438,0.5</points>
<intersection>-4.5 2</intersection>
<intersection>0.5 7</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>454.5,0.5,456.5,0.5</points>
<connection>
<GID>161</GID>
<name>clock</name></connection>
<intersection>454.5 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>438,0.5,438.5,0.5</points>
<connection>
<GID>160</GID>
<name>clock</name></connection>
<intersection>438 5</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>444.5,2.5,444.5,2.5</points>
<connection>
<GID>163</GID>
<name>N_in0</name></connection>
<connection>
<GID>160</GID>
<name>Q</name></connection></vsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>452.5,-1.5,452.5,2.5</points>
<intersection>-1.5 1</intersection>
<intersection>-1.5 1</intersection>
<intersection>2.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>444.5,-1.5,456.5,-1.5</points>
<connection>
<GID>161</GID>
<name>K</name></connection>
<connection>
<GID>160</GID>
<name>nQ</name></connection>
<intersection>452.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>452.5,2.5,456.5,2.5</points>
<connection>
<GID>161</GID>
<name>J</name></connection>
<intersection>452.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>429.5,-27.5,436,-27.5</points>
<connection>
<GID>174</GID>
<name>OUT_0</name></connection>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>432.5 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>432.5,-27.5,432.5,-25</points>
<connection>
<GID>196</GID>
<name>N_in2</name></connection>
<intersection>-27.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>442,-27.5,448.5,-27.5</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<connection>
<GID>176</GID>
<name>OUT_0</name></connection>
<intersection>445 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>445,-27.5,445,-25</points>
<connection>
<GID>198</GID>
<name>N_in2</name></connection>
<intersection>-27.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>454.5,-27.5,462.5,-27.5</points>
<connection>
<GID>178</GID>
<name>OUT_0</name></connection>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>458.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>458.5,-27.5,458.5,-25</points>
<connection>
<GID>200</GID>
<name>N_in2</name></connection>
<intersection>-27.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>423.5,-36,423.5,-30.5</points>
<connection>
<GID>182</GID>
<name>CLK</name></connection>
<connection>
<GID>174</GID>
<name>clock</name></connection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>423.5,-34,462.5,-34</points>
<intersection>423.5 0</intersection>
<intersection>436 6</intersection>
<intersection>448.5 5</intersection>
<intersection>462.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>462.5,-34,462.5,-30.5</points>
<connection>
<GID>180</GID>
<name>clock</name></connection>
<intersection>-34 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>448.5,-34,448.5,-30.5</points>
<connection>
<GID>178</GID>
<name>clock</name></connection>
<intersection>-34 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>436,-34,436,-30.5</points>
<connection>
<GID>176</GID>
<name>clock</name></connection>
<intersection>-34 1</intersection></vsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>423.5,-21,468.5,-21</points>
<intersection>423.5 3</intersection>
<intersection>468.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>423.5,-27.5,423.5,-21</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>-21 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>468.5,-27.5,468.5,-21</points>
<connection>
<GID>180</GID>
<name>OUT_0</name></connection>
<intersection>-23 5</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>468.5,-23,471,-23</points>
<connection>
<GID>206</GID>
<name>N_in0</name></connection>
<intersection>468.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>426.5,-25.5,426.5,-20</points>
<connection>
<GID>174</GID>
<name>set</name></connection>
<connection>
<GID>204</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>430,-59,436.5,-59</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<connection>
<GID>215</GID>
<name>OUT_0</name></connection>
<intersection>433 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>433,-59,433,-56.5</points>
<connection>
<GID>210</GID>
<name>N_in2</name></connection>
<intersection>-59 1</intersection></vsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>442.5,-59,449,-59</points>
<connection>
<GID>217</GID>
<name>IN_0</name></connection>
<connection>
<GID>216</GID>
<name>OUT_0</name></connection>
<intersection>445.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>445.5,-59,445.5,-56.5</points>
<connection>
<GID>211</GID>
<name>N_in2</name></connection>
<intersection>-59 1</intersection></vsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>455,-59,463,-59</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<connection>
<GID>217</GID>
<name>OUT_0</name></connection>
<intersection>459 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>459,-59,459,-56.5</points>
<connection>
<GID>212</GID>
<name>N_in2</name></connection>
<intersection>-59 1</intersection></vsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>424,-67.5,424,-62</points>
<connection>
<GID>219</GID>
<name>CLK</name></connection>
<connection>
<GID>215</GID>
<name>clock</name></connection>
<intersection>-65.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>424,-65.5,463,-65.5</points>
<intersection>424 0</intersection>
<intersection>436.5 6</intersection>
<intersection>449 5</intersection>
<intersection>463 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>463,-65.5,463,-62</points>
<connection>
<GID>218</GID>
<name>clock</name></connection>
<intersection>-65.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>449,-65.5,449,-62</points>
<connection>
<GID>217</GID>
<name>clock</name></connection>
<intersection>-65.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>436.5,-65.5,436.5,-62</points>
<connection>
<GID>216</GID>
<name>clock</name></connection>
<intersection>-65.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>472.5,-59,472.5,-56.5</points>
<connection>
<GID>214</GID>
<name>N_in2</name></connection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>469,-59,472.5,-59</points>
<connection>
<GID>218</GID>
<name>OUT_0</name></connection>
<intersection>472.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>424,-48.5,470.5,-48.5</points>
<intersection>424 4</intersection>
<intersection>470.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>470.5,-62,470.5,-48.5</points>
<intersection>-62 5</intersection>
<intersection>-48.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>424,-59,424,-48.5</points>
<connection>
<GID>215</GID>
<name>IN_0</name></connection>
<intersection>-48.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>469,-62,470.5,-62</points>
<connection>
<GID>218</GID>
<name>OUTINV_0</name></connection>
<intersection>470.5 3</intersection></hsegment></shape></wire></page 4>
<page 5>
<PageViewport>0,126.574,938.642,-337.379</PageViewport></page 5>
<page 6>
<PageViewport>0,126.574,938.642,-337.379</PageViewport></page 6>
<page 7>
<PageViewport>0,126.574,938.642,-337.379</PageViewport></page 7>
<page 8>
<PageViewport>0,126.574,938.642,-337.379</PageViewport></page 8>
<page 9>
<PageViewport>0,126.574,938.642,-337.379</PageViewport></page 9></circuit>